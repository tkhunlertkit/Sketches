module main();

initial
  begin
    $display("Hi there");
    $finish;
  end

endmodule
